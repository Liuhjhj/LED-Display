--	��Ŀ�����޺�Ƶ�·���
--	ʹ��ƽ̨�ϵ�8���߶�����ܽ�����ʾ����Χ��ƽ̨�ϵ�8�������תȦ��
--	Ҫ��ͬʱ��ʾ�Ķ���Ϊ1��2��3�ο�ѡ��
--	�ɽ���˳��������ʾ��ͨ��ĳһ���ؼ�����ѡ�񣩣�
--	���¸�λ�������¿�ʼ��ת��
--	���ֵ�����ʽ��ѡ����ȫ���ȡ�

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LED IS
	PORT(INITLED:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		CLK:IN STD_LOGIC;	--ʱ��ѭ���ź�(��Ƶ��)
		CLR:IN STD_LOGIC;	--��λ�ź�
		FLASH:IN STD_LOGIC;	--ˢ���ź�(��Ƶ��)
		DISPLAY:IN STD_LOGIC_VECTOR(2 DOWNTO 0);	--���ֵ�����ʽѡ��
		ROTATY:IN STD_LOGIC;	--Ϊ1ʱ˳ʱ��,Ϊ0ʱ��ʱ��
		NUMLED:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);	--LED�Ʊ�ţ�0��7
		OUTLED:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));	--LED�ƶ�����0��6
END LED;

ARCHITECTURE DISPLAYLED OF LED IS
SIGNAL COU:INTEGER RANGE 20 DOWNTO 0;
SIGNAL NUM:INTEGER RANGE 0 TO 7;
BEGIN
	PROCESS(FLASH,DISPLAY)	--��Ƶ��
	BEGIN
		IF(DISPLAY/="000" AND DISPLAY/="011" AND DISPLAY/="100" AND DISPLAY/="101") THEN	
			IF(FLASH'EVENT AND FLASH='1') THEN
				IF(NUM=7) THEN
					NUM<=0;
				ELSE
					NUM<=NUM+1;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS(CLK,CLR)	--�޺����ת����Ƶ�ʣ�
	BEGIN
		IF(CLR='1') THEN	--��λ
			COU<=0;
		ELSIF(CLK'EVENT AND CLK='1' AND (DISPLAY="000" OR DISPlAY="011" OR DISPLAY="100" OR DISPLAY="101")) THEN
			IF(COU=20)THEN
				COU<=0;
			ELSE
				COU<=COU+1;
			END IF;
		END IF;
	END PROCESS;
	
	PROCESS(COU)	--�������תȦ
	BEGIN
		IF(DISPLAY="011") THEN	--��ʾ01234567������
			CASE COU IS
				WHEN 0 => NUMLED <= "01111111"; OUTLED <= "1111110";
				WHEN 1 => NUMLED <= "10111111"; OUTLED <= "0110000";
				WHEN 2 => NUMLED <= "11011111"; OUTLED <= "1101101";
				WHEN 3 => NUMLED <= "11101111"; OUTLED <= "1111001";
				WHEN 4 => NUMLED <= "11110111"; OUTLED <= "0110011";
				WHEN 5 => NUMLED <= "11111011"; OUTLED <= "1011011";
				WHEN 6 => NUMLED <= "11111101"; OUTLED <= "1011111";
				WHEN 7 => NUMLED <= "11111110"; OUTLED <= "1110000";
				WHEN OTHERS => NULL;
			END CASE;
		ELSIF(DISPLAY="100") THEN
			NUMLED<="00000000";
			CASE COU IS                                --ѭ����ʾ01234567
				WHEN 0 => OUTLED <= "1111110";
				WHEN 1 => OUTLED <= "0110000";
				WHEN 2 => OUTLED <= "1101101";
				WHEN 3 => OUTLED <= "1111001";
				WHEN 4 => OUTLED <= "0110011";
				WHEN 5 => OUTLED <= "1011011";
				WHEN 6 => OUTLED <= "1011111";
				WHEN 7 => OUTLED <= "1110000";
				WHEN 8 => OUTLED <= "1111111";
				WHEN 9 => OUTLED <= "1111011";
				WHEN OTHERS => OUTLED <= "0000000";
			END CASE;
		ELSIF(DISPLAY="101") THEN						--ѭ����ʾABCDEFGH
			NUMLED<="00000000";
			CASE COU IS
				WHEN 0 => OUTLED <= "1110111";
				WHEN 1 => OUTLED <= "1111111";
				WHEN 2 => OUTLED <= "1001110";
				WHEN 3 => OUTLED <= "1111110";
				WHEN 4 => OUTLED <= "1001111";
				WHEN 5 => OUTLED <= "1000111";
				WHEN 6 => OUTLED <= "1011111";
				WHEN 7 => OUTLED <= "0110111";
				WHEN OTHERS => OUTLED <="0000000";
			END CASE;
			
		ELSIF(DISPLAY="000") THEN
			IF(ROTATY='1') THEN	--˳ʱ����ת
				IF(INITLED="001" OR INITLED="010" OR INITLED="100") THEN	--˳ʱ����һ��
					CASE COU IS
						WHEN 1 => NUMLED <= "01111111"; OUTLED <= "1000000";
						WHEN 2 => NUMLED <= "10111111"; OUTLED <= "1000000";
						WHEN 3 => NUMLED <= "11011111"; OUTLED <= "1000000";
						WHEN 4 => NUMLED <= "11101111"; OUTLED <= "1000000";
						WHEN 5 => NUMLED <= "11110111"; OUTLED <= "1000000";
						WHEN 6 => NUMLED <= "11111011"; OUTLED <= "1000000";
						WHEN 7 => NUMLED <= "11111101"; OUTLED <= "1000000";
						WHEN 8 => NUMLED <= "11111110"; OUTLED <= "1000000";
						WHEN 9 => NUMLED <= "11111110"; OUTLED <= "0100000";
						WHEN 10 =>NUMLED <= "11111110"; OUTLED <= "0010000";
						WHEN 11 =>NUMLED <= "11111110"; OUTLED <= "0001000";
						WHEN 12 =>NUMLED <= "11111101"; OUTLED <= "0001000";
						WHEN 13 =>NUMLED <= "11111011"; OUTLED <= "0001000";
						WHEN 14 =>NUMLED <= "11110111"; OUTLED <= "0001000";
						WHEN 15 =>NUMLED <= "11101111"; OUTLED <= "0001000";
						WHEN 16 =>NUMLED <= "11011111"; OUTLED <= "0001000";
						WHEN 17 =>NUMLED <= "10111111"; OUTLED <= "0001000";
						WHEN 18 =>NUMLED <= "01111111"; OUTLED <= "0001000";
						WHEN 19 =>NUMLED <= "01111111"; OUTLED <= "0000100";
						WHEN 20 =>NUMLED <= "01111111"; OUTLED <= "0000010";
						WHEN  OTHERS => OUTLED <= "0000000";
					END CASE;	
				ELSIF(INITLED="110" OR INITLED="101" OR INITLED="011") THEN	--˳ʱ��������
					CASE COU IS
						WHEN 1 => NUMLED <= "00111111"; OUTLED <= "1000000";
						WHEN 2 => NUMLED <= "11001111"; OUTLED <= "1000000";
						WHEN 3 => NUMLED <= "11110011"; OUTLED <= "1000000";
						WHEN 4 => NUMLED <= "11111100"; OUTLED <= "1000000";
						WHEN 5 => NUMLED <= "11111110"; OUTLED <= "0110000";
						WHEN 6 => NUMLED <= "11111100"; OUTLED <= "0001000";
						WHEN 7 => NUMLED <= "11110011"; OUTLED <= "0001000";
						WHEN 8 => NUMLED <= "11001111"; OUTLED <= "0001000";
						WHEN 9 => NUMLED <= "00111111"; OUTLED <= "0001000";
						WHEN 10=> NUMLED <= "01111111"; OUTLED <= "0000110";
						WHEN OTHERS => OUTLED <= "0000000";
					END CASE;
				ELSIF(INITLED="111") THEN	--˳ʱ��������
					CASE COU IS
						WHEN 1 => NUMLED <= "01111111"; OUTLED <= "1000110";
						WHEN 2 => NUMLED <= "10001111"; OUTLED <= "1000000";
						WHEN 3 => NUMLED <= "11110001"; OUTLED <= "1000000";
						WHEN 4 => NUMLED <= "11111110"; OUTLED <= "1110000";
						WHEN 5 => NUMLED <= "11111000"; OUTLED <= "0001000";
						WHEN 6 => NUMLED <= "11000111"; OUTLED <= "0001000";
						WHEN 7 => NUMLED <= "00111111"; OUTLED <= "0001000";
						WHEN OTHERS => OUTLED <= "0000000";
					END CASE;
				END IF;
			ELSE	--��ʱ����ת
				IF(INITLED="001" OR INITLED="010" OR INITLED="100") THEN	--��ʱ����һ��
					CASE COU IS
						WHEN 20=> NUMLED <= "01111111"; OUTLED <= "1000000";
						WHEN 19=> NUMLED <= "10111111"; OUTLED <= "1000000";
						WHEN 18=> NUMLED <= "11011111"; OUTLED <= "1000000";
						WHEN 17=> NUMLED <= "11101111"; OUTLED <= "1000000";
						WHEN 16=> NUMLED <= "11110111"; OUTLED <= "1000000";
						WHEN 15=> NUMLED <= "11111011"; OUTLED <= "1000000";
						WHEN 14=> NUMLED <= "11111101"; OUTLED <= "1000000";
						WHEN 13=> NUMLED <= "11111110"; OUTLED <= "1000000";
						WHEN 12=> NUMLED <= "11111110"; OUTLED <= "0100000";
						WHEN 11=> NUMLED <= "11111110"; OUTLED <= "0010000";
						WHEN 10=> NUMLED <= "11111110"; OUTLED <= "0001000";
						WHEN 9 => NUMLED <= "11111101"; OUTLED <= "0001000";
						WHEN 8 => NUMLED <= "11111011"; OUTLED <= "0001000";
						WHEN 7 => NUMLED <= "11110111"; OUTLED <= "0001000";
						WHEN 6 => NUMLED <= "11101111"; OUTLED <= "0001000";
						WHEN 5 => NUMLED <= "11011111"; OUTLED <= "0001000";
						WHEN 4 => NUMLED <= "10111111"; OUTLED <= "0001000";
						WHEN 3 => NUMLED <= "01111111"; OUTLED <= "0001000";
						WHEN 2 => NUMLED <= "01111111"; OUTLED <= "0000100";
						WHEN 1 => NUMLED <= "01111111"; OUTLED <= "0000010";
						WHEN  OTHERS => OUTLED <= "0000000";
					END CASE;	
				ELSIF(INITLED="110" OR INITLED="101" OR INITLED="011") THEN	--��ʱ��������
					CASE COU IS
						WHEN 10=> NUMLED <= "00111111"; OUTLED <= "1000000";
						WHEN 9 => NUMLED <= "11001111"; OUTLED <= "1000000";
						WHEN 8 => NUMLED <= "11110011"; OUTLED <= "1000000";
						WHEN 7 => NUMLED <= "11111100"; OUTLED <= "1000000";
						WHEN 6 => NUMLED <= "11111110"; OUTLED <= "0110000";
						WHEN 5 => NUMLED <= "11111100"; OUTLED <= "0001000";
						WHEN 4 => NUMLED <= "11110011"; OUTLED <= "0001000";
						WHEN 3 => NUMLED <= "11001111"; OUTLED <= "0001000";
						WHEN 2 => NUMLED <= "00111111"; OUTLED <= "0001000";
						WHEN 1 => NUMLED <= "01111111"; OUTLED <= "0000110";
						WHEN OTHERS => OUTLED <= "0000000";
					END CASE;
				ELSIF(INITLED="111") THEN	--��ʱ��������
					CASE COU IS
						WHEN 1 => NUMLED <= "01111111"; OUTLED <= "0001110";
						WHEN 2 => NUMLED <= "10001111"; OUTLED <= "0001000";
						WHEN 3 => NUMLED <= "11110001"; OUTLED <= "0001000";
						WHEN 4 => NUMLED <= "11111110"; OUTLED <= "0111000";
						WHEN 5 => NUMLED <= "11111000"; OUTLED <= "1000000";
						WHEN 6 => NUMLED <= "11000111"; OUTLED <= "1000000";
						WHEN 7 => NUMLED <= "00111111"; OUTLED <= "1000000";
						WHEN OTHERS => OUTLED <= "0000000";
					END CASE;
				END IF;
			END IF;
		ELSIF(DISPLAY="001") THEN	--ȫ��
			CASE NUM IS
				WHEN 0 => NUMLED <= "01111111"; OUTLED <= "1001110";
				WHEN 1 => NUMLED <= "10111111"; OUTLED <= "1001000";
				WHEN 2 => NUMLED <= "11011111"; OUTLED <= "1001000";
				WHEN 3 => NUMLED <= "11101111"; OUTLED <= "1001000";
				WHEN 4 => NUMLED <= "11110111"; OUTLED <= "1001000";
				WHEN 5 => NUMLED <= "11111011"; OUTLED <= "1001000";
				WHEN 6 => NUMLED <= "11111101"; OUTLED <= "1001000";
				WHEN 7 => NUMLED <= "11111110"; OUTLED <= "1111000";
				WHEN OTHERS => NULL;
			END CASE;
		ELSIF(DISPLAY="010") THEN	--ͬʱ��ʾ01234567
			CASE NUM IS
				WHEN 0 => NUMLED <= "01111111"; OUTLED <= "1111110";
				WHEN 1 => NUMLED <= "10111111"; OUTLED <= "0110000";
				WHEN 2 => NUMLED <= "11011111"; OUTLED <= "1101101";
				WHEN 3 => NUMLED <= "11101111"; OUTLED <= "1111001";
				WHEN 4 => NUMLED <= "11110111"; OUTLED <= "0110011";
				WHEN 5 => NUMLED <= "11111011"; OUTLED <= "1011011";
				WHEN 6 => NUMLED <= "11111101"; OUTLED <= "1011111";
				WHEN 7 => NUMLED <= "11111110"; OUTLED <= "1110000";
				WHEN OTHERS => NULL;
			END CASE;
		END IF;
	END PROCESS;
	
END ARCHITECTURE DISPLAYLED;

--������:�����������